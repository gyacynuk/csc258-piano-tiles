module VLineRenderer (

);

localparam [8:0] HEIGHT = 9'd480;
localparam [8:0] WIDTH = 9'd240;


endmodule 