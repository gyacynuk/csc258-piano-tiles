module LogicEngine(

);

endmodule 